magic
tech scmos
timestamp 1594499169
<< ntransistor >>
rect -1 16 19 36
<< ndiffusion >>
rect -1 45 19 46
rect -1 37 1 45
rect 7 37 11 45
rect 17 37 19 45
rect -1 36 19 37
rect -1 15 19 16
rect -1 7 1 15
rect 7 7 11 15
rect 17 7 19 15
rect -1 6 19 7
<< ndcontact >>
rect 1 37 7 45
rect 11 37 17 45
rect 1 7 7 15
rect 11 7 17 15
<< polysilicon >>
rect -4 16 -1 36
rect 19 16 22 36
<< metal1 >>
rect -1 37 1 45
rect 7 37 11 45
rect 17 37 19 45
rect -1 7 1 15
rect 7 7 11 15
rect 17 7 19 15
<< end >>
