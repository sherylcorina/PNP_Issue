magic
tech scmos
timestamp 1594543954
<< ntransistor >>
rect -18 192 -8 222
rect -18 142 -8 172
rect -18 92 -8 122
<< ndiffusion >>
rect -18 240 -8 242
rect -18 233 -17 240
rect -10 233 -8 240
rect -18 231 -8 233
rect -18 224 -17 231
rect -10 224 -8 231
rect -18 222 -8 224
rect -18 190 -8 192
rect -18 183 -16 190
rect -9 183 -8 190
rect -18 181 -8 183
rect -18 174 -16 181
rect -9 174 -8 181
rect -18 172 -8 174
rect -18 139 -8 142
rect -18 132 -16 139
rect -9 132 -8 139
rect -18 131 -8 132
rect -18 124 -16 131
rect -9 124 -8 131
rect -18 122 -8 124
rect -18 90 -8 92
rect -18 83 -16 90
rect -9 83 -8 90
rect -18 81 -8 83
rect -18 74 -16 81
rect -9 74 -8 81
rect -18 72 -8 74
<< ndcontact >>
rect -17 233 -10 240
rect -17 224 -10 231
rect -16 183 -9 190
rect -16 174 -9 181
rect -16 132 -9 139
rect -16 124 -9 131
rect -16 83 -9 90
rect -16 74 -9 81
<< polysilicon >>
rect -28 222 -21 228
rect -28 192 -18 222
rect -8 192 -5 222
rect -28 172 -21 178
rect -28 142 -18 172
rect -8 142 -5 172
rect -28 122 -21 128
rect -28 92 -18 122
rect -8 92 -5 122
<< polycontact >>
rect -28 228 -21 235
rect -28 178 -21 185
rect -28 128 -21 135
<< metal1 >>
rect -18 240 -8 241
rect -18 235 -17 240
rect -21 233 -17 235
rect -10 233 -8 240
rect -21 231 -8 233
rect -21 228 -17 231
rect -18 224 -17 228
rect -10 224 -8 231
rect -18 223 -8 224
rect -18 190 -8 191
rect -18 185 -16 190
rect -21 183 -16 185
rect -9 183 -8 190
rect -21 181 -8 183
rect -21 178 -16 181
rect -18 174 -16 178
rect -9 174 -8 181
rect -18 173 -8 174
rect -18 139 -8 141
rect -18 135 -16 139
rect -21 132 -16 135
rect -9 132 -8 139
rect -21 131 -8 132
rect -21 128 -16 131
rect -18 124 -16 128
rect -9 124 -8 131
rect -18 123 -8 124
rect -18 90 -8 91
rect -18 83 -16 90
rect -9 83 -8 90
rect -18 81 -8 83
rect -18 74 -16 81
rect -9 74 -8 81
rect -18 73 -8 74
<< labels >>
rlabel polycontact -23 230 -23 230 3 a
rlabel polycontact -26 182 -26 182 3 b
rlabel polycontact -26 131 -26 131 3 c
<< end >>
