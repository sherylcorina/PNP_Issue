magic
tech scmos
timestamp 1594574876
<< nwell >>
rect -33 -24 27 36
<< pdiffusion >>
rect -13 11 7 16
rect -13 1 -8 11
rect 2 1 7 11
rect -13 -4 7 1
<< pdcontact >>
rect -8 1 2 11
<< psubstratepdiff >>
rect -48 50 42 51
rect -48 42 -47 50
rect -39 42 -32 50
rect -24 42 18 50
rect 26 42 33 50
rect 41 42 42 50
rect -48 41 42 42
rect -48 36 -38 41
rect -48 28 -47 36
rect -39 28 -38 36
rect -48 20 -38 28
rect 32 36 42 41
rect 32 28 33 36
rect 41 28 42 36
rect -48 12 -47 20
rect -39 12 -38 20
rect -48 6 -38 12
rect -48 -2 -47 6
rect -39 -2 -38 6
rect -48 -12 -38 -2
rect -48 -20 -47 -12
rect -39 -20 -38 -12
rect 32 20 42 28
rect 32 12 33 20
rect 41 12 42 20
rect 32 6 42 12
rect 32 -2 33 6
rect 41 -2 42 6
rect 32 -12 42 -2
rect -48 -29 -38 -20
rect 32 -20 33 -12
rect 41 -20 42 -12
rect 32 -29 42 -20
rect -48 -30 42 -29
rect -48 -38 -47 -30
rect -39 -38 -29 -30
rect -21 -38 -12 -30
rect -4 -38 4 -30
rect 12 -38 19 -30
rect 27 -38 33 -30
rect 41 -38 42 -30
rect -48 -39 42 -38
<< nsubstratendiff >>
rect -28 23 -18 26
rect -28 15 -27 23
rect -20 15 -18 23
rect 12 23 22 26
rect -28 8 -18 15
rect -28 0 -27 8
rect -20 0 -18 8
rect -28 -8 -18 0
rect 12 15 14 23
rect 21 15 22 23
rect 12 8 22 15
rect 12 0 14 8
rect 21 0 22 8
rect 12 -8 22 0
rect -28 -9 22 -8
rect -28 -17 -27 -9
rect -20 -17 -17 -9
rect -10 -17 -7 -9
rect 0 -17 4 -9
rect 11 -17 14 -9
rect 21 -17 22 -9
rect -28 -19 22 -17
<< psubstratepcontact >>
rect -47 42 -39 50
rect -32 42 -24 50
rect 18 42 26 50
rect 33 42 41 50
rect -47 28 -39 36
rect 33 28 41 36
rect -47 12 -39 20
rect -47 -2 -39 6
rect -47 -20 -39 -12
rect 33 12 41 20
rect 33 -2 41 6
rect 33 -20 41 -12
rect -47 -38 -39 -30
rect -29 -38 -21 -30
rect -12 -38 -4 -30
rect 4 -38 12 -30
rect 19 -38 27 -30
rect 33 -38 41 -30
<< nsubstratencontact >>
rect -27 15 -20 23
rect -27 0 -20 8
rect 14 15 21 23
rect 14 0 21 8
rect -27 -17 -20 -9
rect -17 -17 -10 -9
rect -7 -17 0 -9
rect 4 -17 11 -9
rect 14 -17 21 -9
<< metal1 >>
rect -39 42 -32 50
rect -47 36 -39 42
rect -47 20 -39 28
rect -47 6 -39 12
rect -47 -12 -39 -2
rect -47 -30 -39 -20
rect -27 23 -20 24
rect -27 8 -20 15
rect -9 11 3 51
rect 26 42 33 50
rect 33 36 41 42
rect -9 1 -8 11
rect 2 1 3 11
rect -9 0 3 1
rect 14 23 21 24
rect 14 8 21 15
rect -27 -9 -20 0
rect 14 -9 21 0
rect -20 -17 -17 -9
rect -10 -17 -7 -9
rect 0 -17 4 -9
rect 11 -17 14 -9
rect -27 -30 21 -17
rect 33 20 41 28
rect 33 6 41 12
rect 33 -12 41 -2
rect 33 -30 41 -20
rect -39 -38 -29 -30
rect -21 -38 -12 -30
rect -4 -38 4 -30
rect 12 -38 19 -30
rect 27 -38 33 -30
<< labels >>
rlabel pdcontact -3 6 -3 6 1 e
rlabel metal1 -2 -18 -2 -18 1 b
<< end >>
